module led(
	output wire [3:0]out		//	4浣嶅淇″彿瀵瑰簲4涓猯ed
);

	assign out[3:0] = 4'b01_01;

	
endmodule